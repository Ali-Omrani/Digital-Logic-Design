module adder(input [15:0]a,b,output [15:0]w);
	assign w=a+b;
	endmodule
	