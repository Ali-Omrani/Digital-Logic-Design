module Q6 (input [15:0] D , N ,output  [15:0] W );
 	
 	assign #(317,289) W = (N[0]==1) ? {D} : 
 	 (N[1]==1) ? {{0},{D[15:1]}} :
 	 (N[2]==1) ? {{2{0}},D[15:2]}:
 	 (N[3]==1) ? {{3{0}},D[15:3]} :
 	 (N[4]==1) ? {{4{0}},D[15:4]} :
 	 (N[5]==1) ? {{5{0}},D[15:5]} :
 	 (N[6]==1) ? {{6{0}},D[15:6]} :
 	 (N[7]==1) ? {{7{0}},D[15:7]} :
 	 (N[8]==1) ? {{8{0}},D[15:8]} :
 	 (N[9]==1) ? {{9{0}},D[15:9]} :
 	 (N[10]==1) ? {{10{0}},D[15:10]} :
 	 (N[11]==1) ? {{11{0}},D[15:11]} :
 	 (N[12]==1) ? {{12{0}},D[15:12]} :
 	 (N[13]==1) ? {{13{0}},D[15:13]} :
 	 (N[14]==1) ? {{14{0}},D[15:14]} :
 	 (N[15]==1) ? {{15{0}},D[15:15]} :0;
 	 
 	 
endmodule