module Q7_testbench();
	logic [15:0] D =16'b1111111111111111;
	logic [15:0] d =1;
	logic [15:0] N =0;
	logic [15:0] n =0;
	logic [15:0] W ;
	logic [15:0] w ;
	
	Q5 MUT1 (D,N,W);	
 	Q6 MUT2 (D,N,w);
	initial begin 
		
		#1000 N[0]=1;
		#1000 N[0]=0;
		N[1]=1;
		#1000 N[1]=0;
		N[2]=1;
		#1000 N[2]=0;
		N[3]=1;
		#1000 N[3]=0;
		N[4]=1;
		#1000 N[4]=0;
		N[5]=1;
		#1000 N[5]=0;
		N[6]=1;
		#1000 N[6]=0;
		N[7]=1;
		#1000 N[7]=0;
		N[8]=1;
		#1000 N[8]=0;
		N[9]=1;
		#1000 N[9]=0;
		N[10]=1;
		#1000 N[10]=0;
		N[11]=1;
		#1000 N[11]=0;
		N[12]=1;
		#1000 N[12]=0;
		N[13]=1;
		#1000 N[13]=0;
		N[14]=1;
		#1000 N[14]=0;
		N[15]=1;
		#1000 N[15]=0;		
		
	end  
endmodule