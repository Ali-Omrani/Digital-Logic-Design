module Q8 (input [7:0] D , N , output [7:0] W);
	nmos #(3,4,5) T1 (W[0],D[0],N[0]);
	nmos #(3,4,5) T2 (W[0],D[1],N[1]);
	nmos #(3,4,5) T3 (W[0],D[2],N[2]);
	nmos #(3,4,5) T4 (W[0],D[3],N[3]);
	nmos #(3,4,5) T5 (W[0],D[4],N[4]);
	nmos #(3,4,5) T6 (W[0],D[5],N[5]);
	nmos #(3,4,5) T7 (W[0],D[6],N[6]);
	nmos #(3,4,5) T8 (W[0],D[7],N[7]);

	nmos #(3,4,5) T9 (W[1],D[7],N[7]);
	nmos #(3,4,5) T10 (W[1],D[1],N[0]);
	nmos #(3,4,5) T11 (W[1],D[2],N[1]);
	nmos #(3,4,5) T12 (W[1],D[3],N[2]);
	nmos #(3,4,5) T13 (W[1],D[4],N[3]);
	nmos #(3,4,5) T14 (W[1],D[5],N[4]);
	nmos #(3,4,5) T15 (W[1],D[6],N[5]);
	nmos #(3,4,5) T16 (W[1],D[7],N[6]);

	nmos #(3,4,5) T17 (W[2],D[7],N[6]);
	nmos #(3,4,5) T18 (W[2],D[7],N[7]);
	nmos #(3,4,5) T19 (W[2],D[2],N[0]);
	nmos #(3,4,5) T20 (W[2],D[3],N[1]);
	nmos #(3,4,5) T21 (W[2],D[4],N[2]);
	nmos #(3,4,5) T22 (W[2],D[5],N[3]);
	nmos #(3,4,5) T23 (W[2],D[6],N[4]);
	nmos #(3,4,5) T24 (W[2],D[7],N[5]);


	nmos #(3,4,5) T25 (W[3],D[7],N[5]);
	nmos #(3,4,5) T26 (W[3],D[7],N[6]);
	nmos #(3,4,5) T27 (W[3],D[7],N[7]);
	nmos #(3,4,5) T28 (W[3],D[3],N[0]);
	nmos #(3,4,5) T29 (W[3],D[4],N[1]);
	nmos #(3,4,5) T30 (W[3],D[5],N[2]);
	nmos #(3,4,5) T31 (W[3],D[6],N[3]);
	nmos #(3,4,5) T32 (W[3],D[7],N[4]);

	nmos #(3,4,5) T33 (W[4],D[7],N[4]);
	nmos #(3,4,5) T34 (W[4],D[7],N[5]);
	nmos #(3,4,5) T35 (W[4],D[7],N[6]);
	nmos #(3,4,5) T36 (W[4],D[7],N[7]);
	nmos #(3,4,5) T37 (W[4],D[4],N[0]);
	nmos #(3,4,5) T38 (W[4],D[5],N[1]);
	nmos #(3,4,5) T39 (W[4],D[6],N[2]);
	nmos #(3,4,5) T40 (W[4],D[7],N[3]);

	nmos #(3,4,5) T41 (W[5],D[7],N[3]);
	nmos #(3,4,5) T42 (W[5],D[7],N[4]);
	nmos #(3,4,5) T43 (W[5],D[7],N[5]);
	nmos #(3,4,5) T44 (W[5],D[7],N[6]);
	nmos #(3,4,5) T45 (W[5],D[7],N[7]);
	nmos #(3,4,5) T46 (W[5],D[5],N[0]);
	nmos #(3,4,5) T47 (W[5],D[6],N[1]);
	nmos #(3,4,5) T48 (W[5],D[7],N[2]);

	nmos #(3,4,5) T49 (W[6],D[7],N[2]);
	nmos #(3,4,5) T50 (W[6],D[7],N[3]);
	nmos #(3,4,5) T51 (W[6],D[7],N[4]);
	nmos #(3,4,5) T52 (W[6],D[7],N[5]);
	nmos #(3,4,5) T53 (W[6],D[7],N[6]);
	nmos #(3,4,5) T54 (W[6],D[7],N[7]);
	nmos #(3,4,5) T55 (W[6],D[6],N[0]);
	nmos #(3,4,5) T56 (W[6],D[7],N[1]);

	nmos #(3,4,5) T57 (W[7],D[7],N[1]);
	nmos #(3,4,5) T58 (W[7],D[7],N[2]);
	nmos #(3,4,5) T59 (W[7],D[7],N[3]);
	nmos #(3,4,5) T60 (W[7],D[7],N[4]);
	nmos #(3,4,5) T61 (W[7],D[7],N[5]);
	nmos #(3,4,5) T62 (W[7],D[7],N[6]);
	nmos #(3,4,5) T63 (W[7],D[7],N[7]);
	nmos #(3,4,5) T64 (W[7],D[7],N[0]);

endmodule